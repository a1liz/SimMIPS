`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/02/2018 08:51:59 AM
// Design Name: 
// Module Name: multiply
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module multiply(
	input wire 			clk,
	input wire 			mult_begin,
	input wire 	[31:0] 	mult_op1,
	input wire 	[31:0] 	mult_op2,
	output wire [63:0] 	product,
	output wire 		mult_end,
	// debug
	output wire         debug_mult_valid,
    output wire [63:0]  debug_product_temp,
    output wire [31:0]  debug_multiplier,
    output wire [31:0]  debug_multiplicand
	);
	
	reg mult_valid;
	assign mult_end = mult_valid & ~(|multiplier);
	always @(posedge clk) 
	begin
		if (!mult_begin || mult_end) 
		begin
			mult_valid <= 1'b0;
		end
		else
		begin
		  mult_valid <= 1'b1;
		end
	end

	wire 		op1_sign;
	wire 		op2_sign;
	wire [31:0] op1_absolute;
	wire [31:0] op2_absolute;
	assign op1_sign = mult_op1[31];
	assign op2_sign = mult_op2[31];
	assign op1_absolute = op1_sign ? (~mult_op1+1) : mult_op1;
    assign op2_absolute = op2_sign ? (~mult_op2+1) : mult_op2;

    //?????????????????????????????????????????????
    reg  [63:0] multiplicand;
    always @ (posedge clk)
    begin
        if (mult_valid)
        begin    // ????????????????????????????????????????????????????????????
            multiplicand <= {multiplicand[62:0],1'b0};
        end
        else if (mult_begin) 
        begin   // ??????????????????????????????????????????1????????????
            multiplicand <= {32'd0,op1_absolute};
        end
    end

    //??????????????????????????????????????????
    reg  [31:0] multiplier;
    always @ (posedge clk)
    begin
        if (mult_valid)
        begin   // ?????????????????????????????????????????????????????????
            multiplier <= {1'b0,multiplier[31:1]}; 
        end
        else if (mult_begin)
        begin   // ???????????????????????????????????????2????????????
            multiplier <= op2_absolute; 
        end
    end
    
    // ???????????????????????????1?????????????????????????????????????????????0???????????????0
    wire [63:0] partial_product;
    assign partial_product = multiplier[0] ? multiplicand : 64'd0;
    
    //?????????
    reg [63:0] product_temp;
    always @ (posedge clk)
    begin
        if (mult_valid)
        begin
            product_temp <= product_temp + partial_product;
        end
        else if (mult_begin) 
        begin
            product_temp <= 64'd0;  // ??????????????????????????? 
        end
    end 
    //???????????????????????????????????????
    reg product_sign;
    always @ (posedge clk)  // ??????
    begin
        if (mult_valid)
        begin
              product_sign <= op1_sign ^ op2_sign;
        end
    end 
    //???????????????????????????????????????????????????+1
    assign product = product_sign ? (~product_temp+1) : product_temp;
    
    // debug
    assign debug_mult_valid = mult_valid;
    assign debug_product_temp = product_temp;
    assign debug_multiplier = multiplier;
    assign debug_multiplicand = multiplicand;
endmodule









